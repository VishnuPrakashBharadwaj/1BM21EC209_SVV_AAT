class transactor;
    function new();
        
    endfunction //new()
endclass //transactor