class receiver;
    task new();
        
    endtask //new()
endclass //receiver