class driver;
    function new();
        
    endfunction //new()
endclass //driver