program counter_test();


endprogram