class receiver;
    function new();
        
    endfunction //new()
endclass //receiver